library IEEE;
use IEEE.std_logic_1164.all;

entity fd is

end entity fd;


architecture rtl of fd is
 
begin
	
	 
end architecture rtl;