library IEEE;
use IEEE.std_logic_1164.all;

entity a is

end entity a;


architecture rtl of a is
 
begin
	
	 
end architecture rtl;